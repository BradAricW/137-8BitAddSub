module su 
(
	input c, p,
	output s
);
	assign s = c ^ p;

endmodule